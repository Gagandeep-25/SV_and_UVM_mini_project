class driver extends uvm_driver#(transaction);
  `uvm_component_utils(driver)
  
  function new(input string path = "driver", uvm_component parent);
    super.new(path,parent);
  endfunction
  
  transaction data;
  virtual add_if aif;
  
  task reset_dut();
    aif.rst <= 1'b1;
    aif.a <= 0;
    aif.b <= 0;
    
    repeat(5) @(posedge aif.clk);
      aif.rst =  1'b0;
    `uvm_info("DRV","Reset Done",UVM_NONE);
  endtask
    
  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    data = transaction::type_id::create("data");
      
    if(!uvm_config_db#(virtual add_if)::get(this,"","aif",aif))
      `uvm_error("DRV","Unable to access");
  endfunction
    
  virtual task run_phase(uvm_phase phase);
    reset_dut();
    forever begin 
      
      seq_item_port.get_next_item(data);
      aif.a <= data.a;
      aif.b <= data.b;
      `uvm_info("DRV",$sformatf("trigger DUT a : %0d and b : %0d",data.a,data.b),UVM_NONE);
      seq_item_port.item_done();
      repeat(2) @(posedge aif.clk); //wait for 2 clk tick unit we send the next transaction to DUT
      
    end
  endtask
  
endclass
