/////////////////////////////////////////////////////////////////////// INTERFACE 
